interface addr_intf(input logic clk,rst);
  
  logic [3:0]a;
  logic [3:0]b;
  logic valid;
  logic [6:0]c;
endinterface
